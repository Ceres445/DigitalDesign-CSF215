`include "demux_1to4"
module full_adder(input [3:0] in,output out);

endmodule
